

`timescale 1ns / 1ps
`default_nettype none


// 以降は Verilator で C++ のテストドライバも使えるように時間待ちを書かない
module tb_main
        (
            input   var logic                       reset   ,
            input   var logic                       clk     
        );


    int     cycle;
    always_ff @( posedge clk ) begin
        if ( reset ) begin
            cycle <= 0;
        end
        else begin
            cycle <= cycle + 1;
            if ( cycle >= 1000 ) begin
                // シミュレーション終了
                automatic int fp = $fopen("simulation_completed.log", "w");
                $fclose(fp);
                $display("Simulation Completed");
                $finish(0);
            end
        end
    end


`ifdef __VERILATOR__
    localparam  DEVICE     = "RTL"              ;   // デバイス名
`else
    localparam  DEVICE     = "ULTRASCALE_PLUS"  ;   // デバイス名
`endif
    localparam  SIMULATION = "true"             ;   // シミュレーション
    localparam  DEBUG      = "false"            ;   // デバッグ


    // -----------------------------------------
    //  SVAを使った parameter別検証
    // -----------------------------------------

    for ( genvar LATENCY = 0; LATENCY <= 3; LATENCY++ ) begin : latency
        for ( genvar N = 2; N <= 32; N++ ) begin : n
            for ( genvar DATA_BITS = 1; DATA_BITS <= 8; DATA_BITS += 8 ) begin : data_bits
                tb_elixirchip_es1_spu_op_sel
                        #(
                            .LATENCY        (LATENCY    ),
                            .N              (N          ),  
                            .DATA_BITS      (DATA_BITS  ),
                            .DEVICE         (DEVICE     ),
                            .SIMULATION     (SIMULATION ),
                            .DEBUG          (DEBUG      )
                        )
                    u_tb_elixirchip_es1_spu_op_sel
                        (
                            .reset          ,
                            .clk            
                        );
            end
        end
    end
    
    // SVA bind  (インスタンスへの bind は verilator が未対応)
    bind elixirchip_es1_spu_op_sel sva_elixirchip_es1_spu_op_sel
            #(
                .LATENCY        (LATENCY    ),
                .DATA_BITS      (DATA_BITS  ),
                .N              (N          ),
                .SEL_BITS       (SEL_BITS   ),
                .CLEAR_DATA     (CLEAR_DATA ),
                .IMMEDIATE_SEL  (1'b0       ),
                .IMMEDIATE_DATA (1'b0       ),
                .DEVICE         (DEVICE     ),
                .SIMULATION     (SIMULATION ),
                .DEBUG          (DEBUG      ) 
            )
        u_sva
            (
                .*
            );


    // -----------------------------------------
    //  typical な個別検証
    // -----------------------------------------

    localparam  int     LATENCY    = 3                       ;   // レイテンシ指定
    localparam  int     N          = 4                       ;   // 入力データ数
    localparam  int     SEL_BITS   = $clog2(N)               ;   // セレクタの幅
    localparam  type    sel_t      = logic [SEL_BITS-1:0]    ;   // データ型指定(オプション)
    localparam  int     DATA_BITS  = 8                       ;   // データ幅指定
    localparam  type    data_t     = logic [DATA_BITS-1:0]   ;   // データ型指定(オプション)
    localparam  data_t  CLEAR_DATA = 123                     ;   // クリア値
    localparam  bit     IMMEDIATE_DATA0 = 1'b0                    ;   // s_data0 が即値の場合に1にする
    localparam  bit     IMMEDIATE_DATA1 = 1'b0                    ;   // s_data1 が即値の場合に1にする

    typedef struct {
        logic           cke     ;   // クロックイネーブル
        sel_t           s_sel   ;   // 選択の入力
        data_t  [N-1:0] s_data  ;   // 入力データ(N個分の配列)
        logic           s_clear ;   // クリア
        logic           s_valid ;   // 信号有効
    } input_signals_t;

    typedef struct {
        data_t          m_data  ;   // 出力データ
    } output_signals_t;

    input_signals_t input_table [] = '{
        '{cke: 1'b1, s_sel: sel_t'(0), s_data: '{8'h03, 8'h02, 8'h01, 8'h00}, s_clear: 1'b0, s_valid: 1'b1}, // 0
        '{cke: 1'b1, s_sel: sel_t'(3), s_data: '{8'h13, 8'h12, 8'h11, 8'h10}, s_clear: 1'b0, s_valid: 1'b1}, // 1
        '{cke: 1'b1, s_sel: sel_t'(1), s_data: '{8'h23, 8'h22, 8'h21, 8'h20}, s_clear: 1'b0, s_valid: 1'b1}, // 2
        '{cke: 1'b1, s_sel: sel_t'(2), s_data: '{8'h33, 8'h32, 8'h31, 8'h30}, s_clear: 1'b0, s_valid: 1'b1}, // 3
        '{cke: 1'b1, s_sel: sel_t'(0), s_data: '{8'h43, 8'h42, 8'h41, 8'h40}, s_clear: 1'b0, s_valid: 1'b1}, // 4
        '{cke: 1'b0, s_sel: sel_t'(1), s_data: '{8'h43, 8'h42, 8'h41, 8'h40}, s_clear: 1'b0, s_valid: 1'b1}, // cke=0 keep
        '{cke: 1'b1, s_sel: sel_t'(1), s_data: '{8'h53, 8'h52, 8'h51, 8'h50}, s_clear: 1'b0, s_valid: 1'b1}, // 5
        '{cke: 1'b1, s_sel: sel_t'(2), s_data: '{8'h63, 8'h62, 8'h61, 8'h60}, s_clear: 1'b0, s_valid: 1'b1}, // 6
        '{cke: 1'b1, s_sel: sel_t'(3), s_data: '{8'h73, 8'h72, 8'h71, 8'h70}, s_clear: 1'b1, s_valid: 1'b1}, // 7 : clear
        '{cke: 1'b1, s_sel: sel_t'(0), s_data: '{8'h83, 8'h82, 8'h81, 8'h80}, s_clear: 1'b0, s_valid: 1'b0}  // 8 : valid=0
    };
    
    output_signals_t expected_table [] = '{
        '{m_data: 8'h00},    // 0
        '{m_data: 8'h13},    // 1
        '{m_data: 8'h21},    // 2
        '{m_data: 8'h32},    // 3
        '{m_data: 8'h40},    // 4
        '{m_data: 8'h51},    // 5
        '{m_data: 8'h62},    // 6
        '{m_data: 8'd123},   // 7
        '{m_data: 8'd123}    // 8
    };

    input_signals_t     in_sig = '{cke: 1'b1, s_sel: sel_t'(0), s_data: '{0, 0, 0, 0}, s_clear: 1'b0, s_valid: 1'b0};
    output_signals_t    out_sig;

    elixirchip_es1_spu_op_sel
            #(
                .LATENCY        (LATENCY    ),
                .N              (N          ),
                .SEL_BITS       (SEL_BITS   ),
                .sel_t          (sel_t      ),
                .DATA_BITS      (DATA_BITS  ),
                .data_t         (data_t     ),
                .CLEAR_DATA     (CLEAR_DATA ),
                .IMMEDIATE_SEL  (1'b0       ),
                .IMMEDIATE_DATA (1'b0       ),
                .DEVICE         (DEVICE     ),
                .SIMULATION     (SIMULATION ),
                .DEBUG          (DEBUG      ) 
            )
        u_elixirchip_es1_spu_op_sel
            (
                .reset      ,
                .clk        ,
                .cke        (in_sig.cke     ),

                .s_sel      (in_sig.s_sel   ),
                .s_data     (in_sig.s_data  ),
                .s_clear    (in_sig.s_clear ),
                .s_valid    (in_sig.s_valid ),

                .m_data     (out_sig.m_data ) 
            );

    int     input_no = 0;
    int     output_no = 0;
    always_ff @( posedge clk ) begin
        if ( reset ) begin
            input_no  <= 0;
            output_no <= -LATENCY - 1;
        end
        else begin
            if ( input_no < input_table.size() ) begin
                in_sig <= input_table[input_no];
            end

            if ( output_no >= 0 &&  output_no < expected_table.size() ) begin
                if ( out_sig.m_data != expected_table[output_no].m_data ) begin
                    $display("ERROR: output_no=%0d m_data=%h expected=%h", output_no, out_sig.m_data, expected_table[output_no].m_data);
                    $finish;
                end
            end
            
            input_no  <= input_no + 1;
            if ( in_sig.cke ) begin
                output_no <= output_no + 1;
                if ( output_no == expected_table.size() - 1 ) begin
                    $display("Single test passed");
                end
            end
        end
    end


endmodule


`default_nettype wire


// end of file
