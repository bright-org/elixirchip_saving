

`timescale 1ns / 1ps
`default_nettype none


// 以降は Verilator で C++ のテストドライバも使えるように時間待ちを書かない
module tb_main
        (
            input   var logic                       reset   ,
            input   var logic                       clk     
        );


    int     cycle;
    always_ff @( posedge clk ) begin
        if ( reset ) begin
            cycle <= 0;
        end
        else begin
            cycle <= cycle + 1;
            if ( cycle >= 3000 ) begin
                // シミュレーション終了
                automatic int fp = $fopen("simulation_completed.log", "w");
                $fclose(fp);
                $display("Simulation Completed");
                $finish(0);
            end
        end
    end

`ifdef __VERILATOR__
    localparam  DEVICE     = "RTL"              ;   // デバイス名
`else
    localparam  DEVICE     = "ULTRASCALE_PLUS"  ;   // デバイス名
`endif
    localparam  SIMULATION = "true"             ;   // シミュレーション
    localparam  DEBUG      = "false"            ;   // デバッグ


    // -----------------------------------------
    //  SVAを使った parameter別検証
    // -----------------------------------------
    
    for ( genvar LATENCY = 0; LATENCY <= 3; LATENCY++ ) begin : latency
        for ( genvar TABLE_SIZE = 2; TABLE_SIZE <= 512; TABLE_SIZE *= 2 ) begin : table_size
            tb_elixirchip_es1_spu_op_lut
                    #(
                        .LATENCY        (LATENCY    ),
                        .TABLE_SIZE     (TABLE_SIZE ),
                        .DATA_BITS      (8          ),
                        .DEVICE         (DEVICE     ),
                        .SIMULATION     (SIMULATION ),
                        .DEBUG          (DEBUG      )
                    )
                u_tb_elixirchip_es1_spu_op_lut
                    (
                        .reset          ,
                        .clk            
                    );
        end
    end
    

    // SVA bind  (インスタンスへの bind は verilator が未対応)
    bind elixirchip_es1_spu_op_lut sva_elixirchip_es1_spu_op_lut
            #(
                .LATENCY        (LATENCY        ),
                .TABLE_SIZE     (TABLE_SIZE     ),
                .ADDR_BITS      (ADDR_BITS      ),
                .DATA_BITS      (DATA_BITS      ),
                .CLEAR_DATA     (CLEAR_DATA     ),
                .TABLE_VALUES   (TABLE_VALUES   ),
                .DEVICE         (DEVICE         ),
                .SIMULATION     (SIMULATION     ),
                .DEBUG          (DEBUG          )
            )
        u_sva
            (
                .*
            );
    

    // -----------------------------------------
    //  typical な個別検証
    // -----------------------------------------

    localparam  int                         LATENCY      = 1                        ;   // レイテンシ指定
    localparam  int                         TABLE_SIZE   = 64                       ;   // テーブルサイズ
    localparam  int                         ADDR_BITS    = $clog2(TABLE_SIZE)       ;   // アドレス幅
    localparam  type                        addr_t       = logic [ADDR_BITS-1:0]    ;   // データ型指定(オプション)
    localparam  int                         DATA_BITS    = 8                        ;   // データ幅指定
    localparam  type                        data_t       = logic [DATA_BITS-1:0]    ;   // データ型指定(オプション)
    localparam  data_t                      CLEAR_DATA   = 123                      ;   // m_data クリア値
    localparam  data_t  [TABLE_SIZE-1:0]    TABLE_VALUES = '{
        8'h00, 8'h01, 8'h02, 8'h03, 8'h04, 8'h05, 8'h06, 8'h07,
        8'h08, 8'h09, 8'h0a, 8'h0b, 8'h0c, 8'h0d, 8'h0e, 8'h0f,
        8'h10, 8'h11, 8'h12, 8'h13, 8'h14, 8'h15, 8'h16, 8'h17,
        8'h18, 8'h19, 8'h1a, 8'h1b, 8'h1c, 8'h1d, 8'h1e, 8'h1f,
        8'h20, 8'h21, 8'h22, 8'h23, 8'h24, 8'h25, 8'h26, 8'h27,
        8'h28, 8'h29, 8'h2a, 8'h2b, 8'h2c, 8'h2d, 8'h2e, 8'h2f,
        8'h30, 8'h31, 8'h32, 8'h33, 8'h34, 8'h35, 8'h36, 8'h37,
        8'h38, 8'h39, 8'h3a, 8'h3b, 8'h3c, 8'h3d, 8'h3e, 8'h3f
    };

    typedef struct {
        logic   cke     ;   // クロックイネーブル
        addr_t  s_addr  ;   // キャリー入力
        logic   s_clear ;   // クリア
        logic   s_valid ;   // 信号有効
    } input_signals_t;

    typedef struct {
        data_t  m_data  ;   // 出力データ
    } output_signals_t;

    input_signals_t input_table [] = '{
        '{cke: 1'b1, s_addr: addr_t'(   0), s_clear: 1'b0, s_valid: 1'b1},    // 0 
        '{cke: 1'b1, s_addr: addr_t'(  63), s_clear: 1'b0, s_valid: 1'b1},    // 1 
        '{cke: 1'b1, s_addr: addr_t'(   1), s_clear: 1'b0, s_valid: 1'b1},    // 2 
        '{cke: 1'b1, s_addr: addr_t'(   2), s_clear: 1'b1, s_valid: 1'b1},    // 3 clear
        '{cke: 1'b1, s_addr: addr_t'(   3), s_clear: 1'b0, s_valid: 1'b1},    // 4 
        '{cke: 1'b0, s_addr: addr_t'(   4), s_clear: 1'b0, s_valid: 1'b1},    // cke=0 keep
        '{cke: 1'b1, s_addr: addr_t'(   5), s_clear: 1'b0, s_valid: 1'b0},    // 5 valid=0
        '{cke: 1'b1, s_addr: addr_t'(   6), s_clear: 1'b0, s_valid: 1'b1}     // 6 
    };
    
    output_signals_t expected_table [] = '{
        '{m_data: data_t'(63 -  0)},  // 0
        '{m_data: data_t'(63 - 63)},  // 1
        '{m_data: data_t'(63 -  1)},  // 2
        '{m_data: data_t'(    123)},  // 3
        '{m_data: data_t'(63 -  3)},  // 4
        '{m_data: data_t'(63 -  3)},  // 5
        '{m_data: data_t'(63 -  6)}   // 6
    };

    input_signals_t     in_sig = '{cke: 1'b1, s_addr: addr_t'(0), s_clear: 1'b0, s_valid: 1'b0};
    output_signals_t    out_sig;

    elixirchip_es1_spu_op_lut
            #(
                .LATENCY        (LATENCY        ),
                .TABLE_SIZE     (TABLE_SIZE     ),
                .ADDR_BITS      (ADDR_BITS      ),
                .addr_t         (addr_t         ),
                .DATA_BITS      (DATA_BITS      ),
                .data_t         (data_t         ),
                .CLEAR_DATA     (CLEAR_DATA     ),
                .TABLE_VALUES   (TABLE_VALUES   ),
                .USE_CLEAR      (1'b1           ),
                .USE_VALID      (1'b1           ),
                .DEVICE         (DEVICE         ),
                .SIMULATION     (SIMULATION     ),
                .DEBUG          (DEBUG          )
            )
        u_elixirchip_es1_spu_op_lut
            (
                .reset   ,
                .clk     ,
                .cke     (in_sig.cke      ),

                .s_addr  (in_sig.s_addr   ),
                .s_clear (in_sig.s_clear  ),
                .s_valid (in_sig.s_valid  ),

                .m_data  (out_sig.m_data  ) 
            );

    int     input_no = 0;
    int     output_no = 0;
    always_ff @( posedge clk ) begin
        if ( reset ) begin
            input_no  <= 0;
            output_no <= -LATENCY - 1;
        end
        else begin
            if ( input_no < input_table.size() ) begin
                in_sig <= input_table[input_no];
            end

            if ( output_no >= 0 &&  output_no < expected_table.size() ) begin
                if ( out_sig.m_data != expected_table[output_no].m_data ) begin
                    $display("ERROR: output_no=%0d m_data=%h expected=%h", output_no, out_sig.m_data, expected_table[output_no].m_data);
                    $finish;
                end
            end
            
            input_no  <= input_no + 1;
            if ( in_sig.cke ) begin
                output_no <= output_no + 1;
                if ( output_no == expected_table.size() - 1 ) begin
                    $display("Single test passed");
                end
            end
        end
    end

endmodule


`default_nettype wire


// end of file
